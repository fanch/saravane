msgid ""
msgstr ""
"Project-Id-Version: NuTyX Configuration tool\n"
"PO-Revision-Date: 2014-08-07+2000\n"
"Last-Translator: https://translate.google.se/#fr/sv/\n"
"Language-Team: Swedish\n"
"Language: sv \n"
"MIME-Version: 1.0\n"
"Content-Type: text/plain; charset=UTF-8\n"
"Content-Transfer-Encoding: 8bit\n"

msgid "Settings"
msgstr "Inställningar"

msgid "Keyboard Layout"
msgstr "Tangentbordslayout"

msgid "Choose available"
msgstr "Välj tillgängliga"

msgid "ERROR configuration"
msgstr "ERROR konfiguration"

msgid "Please try again"
msgstr "Försök igen"

msgid "Network card"
msgstr "Nätverkskort"

msgid "Select the card"
msgstr "Välj det kort"

msgid "Card to configure"
msgstr "Kort för att konfigurera"

msgid "Configuration of"
msgstr "Konfiguration av"

msgid "Configuration mode"
msgstr "Konfigurationsläge"

msgid "Auto"
msgstr "Auto"

msgid "Man"
msgstr "Man"

msgid "IP address automatically set from DHCP server"
msgstr "IP adress automatiskt från DHCP-servern"

msgid "Manually specify parameters"
msgstr "Ange parametrar manuellt"

msgid "Enter an IP address"
msgstr "Ange en IP-adress"

msgid "Enter a broadcast address"
msgstr "Ange en broadcast-adress"

msgid "in most cases the current value can be used"
msgstr "i de flesta fall det aktuella värdet kan användas"

msgid "Enter the subnet mask"
msgstr "Ange nätmasken"

msgid "Enter the gateway address"
msgstr "Ange gateway-adress"

msgid "it is normally the address of your router access point"
msgstr "Det är normalt den adressen för din router åtkomstpunkt"

msgid "Enter the DNS address"
msgstr "Ange DNS-adress"

msgid "DNS Search Suffix"
msgstr "DNS-sökning Suffix"

msgid "Enter the domain name"
msgstr "Ange det domännamn"

msgid "this is only need if you are in a subdomain"
msgstr "detta behöver bara om du är i en underdomän"

msgid "Most of the time it's not need"
msgstr "Merparten av tiden det inte behöver"

msgid "Start the service"
msgstr "Starta tjänsten"

msgid "Check the all configuration, return true or false"
msgstr "Kontrollera all konfiguration, returnera sant eller falskt"

msgid "Show the network configuration"
msgstr "Visa nätverkskonfigurationen"

msgid "Show the keyboard configuration"
msgstr "Visa tangentbordskonfigurationen"

msgid "Show the clock configuration"
msgstr "Visar konfigurationen klockan"

msgid "Show the locale and local time adjustment"
msgstr "Visa lokalen och lokal tid justering"

msgid "Show the all configuration"
msgstr "Visar all konfiguration"

msgid "Configure the language"
msgstr "Konfigurerar språket"

msgid "Configure the keyboard"
msgstr "Konfigurera tangentbordet"

msgid "Configure the network"
msgstr "Konfigurera nätverket"

msgid "Configure the clock"
msgstr "Konfigurera klocka"

msgid "add a user to the system"
msgstr "lägga till en användare i systemet"

msgid "Configure the all system"
msgstr "Konfigurera all system"

msgid "Install NuTyX"
msgstr "Installera NuTyX"

msgid "Use the arrows keys to change the values"
msgstr "Använd piltangenterna för att ändra värdena"

msgid "Coordinated Universal Time or Local Time ?"
msgstr "Coordinated Universal Time eller Lokal tid ?"

msgid "The hardware clock is set to"
msgstr "Maskinvaruklockan är inställd på"

msgid "Do you want to use this time as Coordinated Universal Time ?"
msgstr "Vill du använda denna tid som Coordinated Universal Time ?"

msgid "and have the summer/winter time changing automatically"
msgstr "och har sommar / vintertid förändras automatiskt"

msgid "Please enter the date"
msgstr "Vänligen ange datum"

msgid "Please enter the time"
msgstr "Ange tiden"

msgid "Configuration of the boot of the machine (GRUB)"
msgstr "Konfiguration av bagageutrymmet på maskinen (GRUB)"

msgid "Select the disk on which you want to modify the MBR"
msgstr "Välj den disk som du vill ändra MBR"

msgid "Select the partition on which should be located the GRUB files"
msgstr "Välj den partition som ska placeras på GRUB-filer"

msgid "Note that the destination partition can contain NuTyX or any other distribution"
msgstr "Observera att destinationen partition kan innehålla NuTyX eller någon annan distribution"

msgid "No boot process configured"
msgstr "Ingen startprocessen konfigureras"

msgid "You have installed NuTyX without configuring the boot process"
msgstr "Du har installerat NuTyX utan konfiguration av startprocessen"

msgid "Are you sure, you want to cancel the process ?"
msgstr "Är du säker på att du vill avbryta processen ?"

msgid "You already have a copy of the original MBR, it will not be backup"
msgstr "Du har redan en kopia av den ursprungliga MBR, kommer det inte vara backup"

msgid "Good to know"
msgstr "Bra att veta"

msgid "Main Menu"
msgstr "Huvudmeny"

msgid "Welcome in the NuTyX installer"
msgstr "Välkommen i NuTyX installations"

msgid "Create all your partitions"
msgstr "Skapa alla dina partition"

msgid "Format a partition"
msgstr "Formatera en partition"

msgid "Configure the boot of the PC"
msgstr "Konfigurera bagageutrymmet på datorn"

msgid "Reboot the PC"
msgstr "Starta om datorn"

